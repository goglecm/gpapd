library ieee;
use ieee.std_logic_1164.all;

---------------------------------------

entity c_element is
    port
    (
        a_in  : in  std_ulogic;
        b_in  : in  std_ulogic;
        c_out : out std_ulogic
    );
end entity;
